module  SMS_CARD_HIZ(
    output a 
    );

    assign a = 1'bz;

endmodule

module  SMS_CARD_ONE(
    output a 
    );

    assign a = 1;

endmodule

module  SMS_CARD_ZERO(
    output a 
    );

    assign a = 0;

endmodule
